
  `ifndef _MAIN_PARAMETERS_
  `define _MAIN_PARAMETERS_

  `define _FREQ_CLK_        50000000
  `define _LEDS_WIDTH_      8
  `define _BUTTONS_WIDTH_   2
  `define _SWITCHES_WIDTH_  4
  `define _GPIO_0_WIDTH_    36
  `define _GPIO_1_WIDTH_    36

  `endif
