
  `ifndef _AXI_SPI_DEFINES_
  `define _AXI_SPI_DEFINES_

  `define _AXI_SPI_DATA_WIDTH_  32
  `define _AXI_SPI_ADDR_WIDTH_  7
  `define _AXI_SPI_FIFO_DEPTH_  32
  `define _AXI_SPI_RESP_WIDTH_  2
  `define _AXI_SPI_ID_WIDTH_    12

  `endif
